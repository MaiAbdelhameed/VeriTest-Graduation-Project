module simple_not (
  input in,
  output out
);

  assign out = ~in; // Invert the input

endmodule