module not8 (
  input in,
  output out
);

  nor (out, in, in);

endmodule