module and6 (
    input wire a,
    output wire out
);

assign out = (a == 1'b1);

endmodule
