module parameterized_state_machine #(parameter IDLE = 3'b000, ACTIVE = 3'b001, DONE = 3'b010) (
  // ... same structure as previous examples, using IDLE, ACTIVE, DONE in case statements
);
