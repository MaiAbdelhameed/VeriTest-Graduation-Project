// tested
module and1 (
  input a,
  input b,
  output out
);

  assign out = a & b; // Performs an AND operation

endmodule
