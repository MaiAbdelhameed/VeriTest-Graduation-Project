module simple_and (
  input a,
  input b,
  output out
);

  assign out = a & b; // Performs an AND operation

endmodule
