// tested
module or2_gate (
  input a,
  input b,
  output out
);

  // Instantiate an OR gate primitive
  or (out, a, b);

endmodule