module not5 (
  input in,
  output out
);

  nand (out, in, in);

endmodule