// tested
module and14 (
    input wire [2:0] a,
    input wire [2:0] b,
    output reg [2:0] out
);
    always @(*) begin
        out = {a[2] & b[2], a[1] & b[1], a[0] & b[0]};
    end

endmodule
