//built-in operator
module simple_or (
  input a,
  input b,
  output out
);

  assign out = a | b;

endmodule