module simple_xor (
  input a,
  input b,
  output out
);

  assign out = a ^ b; // ^ represents the XOR operator

endmodule