// tested
module and12 (
    input wire [3:0] a,
    input wire [3:0] b,
    output wire [3:0] out
);

integer i;

always @(*) begin
    for (i = 0; i < 4; i = i + 1) begin
        out[i] = a[i] & b[i];
    end
end


endmodule
