module gate_not (
  input in,
  output out
);

  not (out, in); // Instantiate a NOT gate primitive

endmodule