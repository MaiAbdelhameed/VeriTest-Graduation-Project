// 6 input and
// tested
module and23 (
  input a,
  input b,
  input c,
  input d,
  input e,
  input f,
  output out
);

  assign out = a & b & c & d & e & f; // Performs an AND operation

endmodule
