// 8 input and
// tested
module and30 (
  input a,
  input b,
  input c,
  input d,
  input e,
  input f,
  input g,
  input h,
  output out
);

  assign out = &{a,b,c,d,e,f,g,h}; // Performs an AND operation

endmodule
