module unary_and_bitwise(
    input wire a,
    output wire out
);

assign out = &a;

endmodule
