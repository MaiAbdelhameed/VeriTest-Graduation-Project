module mult10 (input a, b,
            output result); // tested

    assign result = a&b;
endmodule