module mult14(input a, b,
            output result);

    assign result = a&b;
endmodule